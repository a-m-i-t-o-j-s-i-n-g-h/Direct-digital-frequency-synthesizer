module LUT_ROM #(
    parameter n = 18,
    parameter l = 6
)(
    input  wire [l-1:0] phi_lut,    
    input  wire       LM,          
    output wire [63:0] lut_data   
);

    wire [3:0] addr_lut0 = phi_lut[l-1 -: 4]; 
    wire [5:0] addr_lut1 = phi_lut;      

    reg [63:0] ROM0 [0:15];  
    reg [63:0] ROM1 [0:63];  

    reg [63:0] data_out;

    initial begin
        ROM0[ 0] = 64'h8000000000648000;
        ROM0[ 1] = 64'h7FD3106B2F646054;
        ROM0[ 2] = 64'h7F4C80D6136400A8;
        ROM0[ 3] = 64'h7E6C9140616350FC;
        ROM0[ 4] = 64'h7D33F1A9CE62514E;
        ROM0[ 5] = 64'h7BA37212106121A0;
        ROM0[ 6] = 64'h79BC4278DE5FA1F1;
        ROM0[ 7] = 64'h777F92DDF05DE240;
        ROM0[ 8] = 64'h74EF1340FF5BD28E;
        ROM0[ 9] = 64'h720C83A1C65992DA;
        ROM0[10] = 64'h6ED9F40000571324;
        ROM0[11] = 64'h6B59945B6C54536C;
        ROM0[12] = 64'h678DE4B3C95153B1;
        ROM0[13] = 64'h63798508D94E23F4;
        ROM0[14] = 64'h5F1F655A614AB434;
        ROM0[15] = 64'h5A8285A828471471;


    end

    initial begin
ROM1[0]  = 64'h8000000000648000;
ROM1[1]  = 64'h7FFD701988648014;
ROM1[2]  = 64'h7FF5D0330F648028;
ROM1[3]  = 64'h7FE9104C9464703C;
ROM1[4]  = 64'h7FD7406616646050;
ROM1[5]  = 64'h7FC0607F93645064;
ROM1[6]  = 64'h7FA460990C644078;
ROM1[7]  = 64'h7F8350B27F64208C;
ROM1[8]  = 64'h7F5D30CBEA6410A0;
ROM1[9]  = 64'h7F31F0E54E63E0B4;
ROM1[10] = 64'h7F01B0FEA863C0C8;
ROM1[11] = 64'h7ECC6117F86390DC;
ROM1[12] = 64'h7E9201313D6370F0;
ROM1[13] = 64'h7E52A14A76633104;
ROM1[14] = 64'h7E0E3163A2630117;
ROM1[15] = 64'h7DC4C17CBF62C12B;
ROM1[16] = 64'h7D765195CE62913F;
ROM1[17] = 64'h7D22E1AECC625152;
ROM1[18] = 64'h7CCA71C7B9620166;
ROM1[19] = 64'h7C6D11E09461C179;
ROM1[20] = 64'h7C0AC1F95C61718D;
ROM1[21] = 64'h7BA37212106121A0;
ROM1[22] = 64'h7B37422AAE60C1B4;
ROM1[23] = 64'h7AC63243376071C7;
ROM1[24] = 64'h7A50325BA96D11DA;
ROM1[25] = 64'h79D56274025FB1ED;
ROM1[26] = 64'h7955B28C435F5200;
ROM1[27] = 64'h78D132A4695EE213;
ROM1[28] = 64'h7847E2BC755E7226;
ROM1[29] = 64'h77B9C2D4655E1239;
ROM1[30] = 64'h7726E2EC385D924C;
ROM1[31] = 64'h768F4303ED5D225E;
ROM1[32] = 64'h75F2F31B845CA271;
ROM1[33] = 64'h7551F332FB5C2283;
ROM1[34] = 64'h74AC434A515BA296;
ROM1[35] = 64'h7401E361865B22A8;
ROM1[36] = 64'h7352F378985A92BA;
ROM1[37] = 64'h729F738F875A02CC;
ROM1[38] = 64'h71E753A6525972DE;
ROM1[39] = 64'h712AB3BCF758E2F0;
ROM1[40] = 64'h706993D377585301;
ROM1[41] = 64'h6FA3F3E9CF57B313;
ROM1[42] = 64'h6ED9F40000571324;
ROM1[43] = 64'h6E0B741608567336;
ROM1[44] = 64'h6D38A42BE655D347;
ROM1[45] = 64'h6C6174419A552358;
ROM1[46] = 64'h6B86045722547369;
ROM1[47] = 64'h6AA6346C7F53C379;
ROM1[48] = 64'h69C23481AE53138A;
ROM1[49] = 64'h68DA0496AF52639B;
ROM1[50] = 64'h67ED94AB8251A3AB;
ROM1[51] = 64'h66FD14C02550E3BB;
ROM1[52] = 64'h660874D4975023CB;
ROM1[53] = 64'h650FC4E8D94F63DB;
ROM1[54] = 64'h641314FCE84EA3EB;
ROM1[55] = 64'h63126510C54DD3FA;
ROM1[56] = 64'h620DC5246E4D040A;
ROM1[57] = 64'h61053537E24C3419;
ROM1[58] = 64'h5FF8D54B224B6428;
ROM1[59] = 64'h5EE8A55E2C4A9437;
ROM1[60] = 64'h5DD4A570FE49B446;
ROM1[61] = 64'h5CBCF5839A48D455;
ROM1[62] = 64'h5BA18595FD47F463;
ROM1[63] = 64'h5A8285A828471471;
    end

    always @(*) begin
        case (LM)
            1'b0: data_out = ROM0[addr_lut0];
            1'b1: data_out = ROM1[addr_lut1];
            default: data_out = 64'b0;
        endcase
    end

    assign lut_data = data_out;

endmodule
